module IF_ID_reg();

endmodule